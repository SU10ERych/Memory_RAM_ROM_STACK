
`timescale 1ns/1ns
module testbench;

	reg [15:0] data_in;
	reg [7:0] addr;
	reg we;
	reg clk;
	reg byteena;
	wire [15:0] data_out;
	wire [7:0] addr_out;

	RAM dut (data_in, addr, we, clk, byteena, data_out, addr_out);
	initial
		begin
			byteena = 0;
			clk = 0;
			we = 0;
			addr = 8'b00000000;
			data_in = 16'b0000000000000000;

			#40; we = 0; byteena = 0;
			for (addr=0; addr < 8; addr= addr+1)
				begin
					#40;
					data_in = data_in + 16'b0010000000000000;
				end

			#40; we = 0; byteena = 1; data_in = 16'b0000000000000000;
			for (addr=0; addr < 8; addr= addr+1)
				begin
					#40;
					data_in = data_in + 16'b0000100000000000;
				end
				#40;
		end

		always #10 clk = ~clk;
		initial
			#600 $finish;

		initial
			$monitor("data_in=%b addr=%b we=%b clk=%b data_out=%b addr_out=%b", data_in, addr, we, clk, data_out, addr_out);
 
		initial
			$dumpvars;
endmodule
